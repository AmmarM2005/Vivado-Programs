module or_gate_gatelevel(input A,B, output Z);
or(Z,A,B);
endmodule