module and_gate_Gatelevel(input A,B,output Z);
and(Z,A,B);
endmodule